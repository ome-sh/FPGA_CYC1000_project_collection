
module clk (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
